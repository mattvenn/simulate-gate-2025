Standard cell Simulation
* this file edited to remove everything not in tt lib
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* include the standard cells
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

* instantiate the cell - adjust this to match your standard cell
Xcell A B VGND VGND VPWR VPWR Y sky130_fd_sc_hd__nand2_1

* use an inverter as a load for the cell to drive
Xnot  Y VGND VGND VPWR VPWR NOTY sky130_fd_sc_hd__inv_1

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse for A and B
* parameters are: initial value, pulsed value, delay time, rise time, fall time, pulse width, period
Va A VGND pulse(0 1.8 1n   10p 10p 1n 2n)
Vb B VGND pulse(0 1.8 1.5n 10p 10p 1n 2n)

* setup the transient analysis
.tran 10p 3n 0

.control
run
set color0 = white
set color1 = black
plot A B Y
.endc

.end
