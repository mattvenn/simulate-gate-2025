Standard cell Simulation
* this file edited to remove everything not in tt lib
.lib "/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* include the standard cells
.include /foss/pdks/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

* instantiate the cell - adjust this to match your standard cell
Xcell A B VGND VGND VPWR VPWR Y sky130_fd_sc_hd__nand2_1

* set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

* create pulse for A and B
* parameters are: initial value, pulsed value, delay time, rise time, fall time, pulse width, period
Va A VGND pulse(0 1.8 1n   10p 10p 1n 2n)
Vb B VGND pulse(0 1.8 1.5n 10p 10p 1n 2n)

* setup the transient analysis
.tran 10p 3n 0

.control
run

set color0 = white
set color1 = black
set color1 = green
set hcopypscolor        ; enable color in PostScript
set hcopydevtype = svg
hardcopy nand.svg A B Y

meas tran y0 AVG y from=0.2n to=0.4n > check.txt
meas tran y1 AVG y from=0.6n to=0.8n >> check.txt
meas tran y2 AVG y from=1.2n to=1.4n >> check.txt
meas tran y3 AVG y from=1.6n to=1.8n >> check.txt
meas tran y4 AVG y from=2.2n to=2.4n >> check.txt
meas tran y5 AVG y from=2.6n to=2.8n >> check.txt

quit
.endc

.end
